package slv_pkg;
//  `include "stimulator.sv"
//  `include "monitor.sv"
//  `include "checker.sv"
//  `include "env.sv"

class stimulator;
endclass

class monitor;
endclass

class chker;
endclass

class env;
endclass
endpackage
