

package fmt_pkg;
  `include "fmt_ini_trans.sv"
  `include "fmt_rsp_trans.sv"
  `include "fmt_ini_mon.sv"
  `include "fmt_rsp_mon.sv"
  //`include "fmt_checker.sv"
  `include "fmt_checker2.sv"
endpackage
