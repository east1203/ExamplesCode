
class slv_trans;
  logic [31:0] data;
endclass
