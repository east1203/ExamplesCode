
package rpt_pkg;
  import report_pkg::*;

  `include "rpt_stm.sv"
  `include "rpt_mon.sv"
  `include "rpt_checker.sv"
  `include "rpt_env.sv"
endpackage
