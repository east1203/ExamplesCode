
package slv_pkg;
  `include "slv_trans.sv"
  `include "slv_ini_mon.sv"
  `include "slv_rsp_mon.sv"
endpackage
